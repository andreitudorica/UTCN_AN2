[aimspice]
[description]
453
NAND with bipolar

.MODEL TRANS NPN TR=5e-9 TF=8e-9
.MODEL DIODE D TT=5e-9 

VCC VCC 0 DC 5

*AC MODE
*VA A 0 PULSE(0.1 4.9 0 1e-10 1e-10 1e-7 2e-7)
*VB B 0 PULSE(0.2 4.8 0 1e-10 1e-10 2e-7 4e-7)

*DC MODE
VA A 0 DC 5
VB B 0 DC 5


D1 0 A DIODE
D2 0 B DIODE

Q11 2 1 A TRANS
Q12 2 1 B TRANS
R1 VCC 1 4k

R2 VCC 3 1.6k
Q2 3 2 4 TRANS
R4 4 0 1k

R3 VCC 5 130
Q3 5 3 6 TRANS
D3 6 OUT DIODE
Q4 OUT 4 0 TRANS

COUT OUT 0 15p

[dc]
1
VA
0
5
0.1
[tran]
1e-9
7e-7
X
X
0
[ana]
1 2
0
1 1
1 1 0 5
4
v(2)
v(3)
v(4)
v(out)
0
1 1
1 1 -0.03 0
1
i(vcc)
[end]
